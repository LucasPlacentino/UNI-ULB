** Profile: "SCHEMATIC1-BIAS"  [ C:\Users\lucasp\repo\UNI-ULB\BA3\ELEC-H314\labo\Labo1\Labo 1 source commune\ampli source commune-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "BIAS.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/lucasp/repo/UNI-ULB/BA3/ELEC-H314/labo/Labo1/libraries for elec-h402/ald.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
